module OR(out1,in1,in2); 
input in1,in2; 
output logic out1; 

assign out1 = in1 | in2; 

endmodule 